CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 110 6 70 10
177 88 765 812
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
345 184 458 281
9437202 0
0
6 Title:
5 Name:
0
0
0
10
6 74LS48
188 796 207 0 14 29
0 3 6 5 4 17 18 8 9 10
11 12 13 14 19
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 976 274 0 18 19
10 14 13 12 11 10 9 8 20 21
1 1 1 1 1 1 1 2 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9998 0 0
2
43530.4 1
0
9 2-In AND~
219 621 160 0 3 22
0 7 6 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3536 0 0
2
43530.4 2
0
9 2-In AND~
219 451 167 0 3 22
0 4 5 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4597 0 0
2
43530.4 3
0
2 +V
167 258 167 0 1 3
0 2
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
43530.4 4
0
7 Pulser~
4 161 266 0 10 12
0 22 23 24 15 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
5.89883e-315 0
0
6 74112~
219 704 277 0 7 32
0 2 16 15 16 2 25 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5616 0 0
2
5.89883e-315 5.26354e-315
0
6 74112~
219 542 277 0 7 32
0 2 7 15 7 2 26 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9323 0 0
2
5.89883e-315 5.30499e-315
0
6 74112~
219 400 277 0 7 32
0 2 4 15 4 2 27 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
317 0 0
2
5.89883e-315 5.32571e-315
0
6 74112~
219 239 277 0 7 32
0 2 28 15 29 2 30 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3108 0 0
2
5.89883e-315 5.34643e-315
0
35
7 7 0 0 0 0 0 1 2 0 0 5
828 171
1018 171
1018 333
991 333
991 310
8 6 0 0 0 0 0 1 2 0 0 5
828 180
1013 180
1013 328
985 328
985 310
9 5 0 0 0 0 0 1 2 0 0 5
828 189
1008 189
1008 323
979 323
979 310
10 4 0 0 0 0 0 1 2 0 0 5
828 198
930 198
930 338
973 338
973 310
11 3 0 0 0 0 0 1 2 0 0 5
828 207
935 207
935 333
967 333
967 310
12 2 0 0 0 0 0 1 2 0 0 5
828 216
940 216
940 328
961 328
961 310
13 1 0 0 0 0 0 1 2 0 0 5
828 225
945 225
945 323
955 323
955 310
1 0 2 0 0 4096 0 9 0 0 22 2
400 214
400 205
7 1 3 0 0 8320 0 7 1 0 0 4
728 241
753 241
753 171
764 171
0 4 4 0 0 8320 0 0 1 25 0 3
330 241
330 198
764 198
0 3 5 0 0 12416 0 0 1 32 0 4
426 240
440 240
440 189
764 189
0 2 6 0 0 12416 0 0 1 31 0 4
590 241
621 241
621 180
764 180
0 0 2 0 0 4096 0 0 0 16 22 2
633 289
633 205
0 0 2 0 0 0 0 0 0 17 22 2
451 289
451 205
0 0 2 0 0 0 0 0 0 22 18 2
312 205
312 289
5 5 2 0 0 4096 0 8 7 0 0 2
542 289
704 289
5 5 2 0 0 4096 0 9 8 0 0 2
400 289
542 289
5 5 2 0 0 4096 0 10 9 0 0 2
239 289
400 289
2 0 7 0 0 4096 0 8 0 0 20 2
518 241
505 241
4 3 7 0 0 16512 0 8 4 0 0 5
518 259
505 259
505 241
472 241
472 167
1 0 2 0 0 16 0 8 0 0 22 2
542 214
542 205
1 0 2 0 0 8320 0 7 0 0 23 3
704 214
704 205
258 205
1 1 2 0 0 0 0 10 5 0 0 4
239 214
239 205
258 205
258 176
2 0 4 0 0 0 0 9 0 0 25 2
376 241
355 241
7 0 4 0 0 0 0 10 0 0 26 2
263 241
355 241
1 4 4 0 0 0 0 4 9 0 0 4
427 158
355 158
355 259
376 259
3 0 15 0 0 8192 0 10 0 0 35 3
209 250
208 250
208 302
3 1 7 0 0 0 0 4 3 0 0 3
472 167
472 151
597 151
2 0 16 0 0 4096 0 7 0 0 30 2
680 241
653 241
3 4 16 0 0 8320 0 3 7 0 0 4
642 160
653 160
653 259
680 259
7 2 6 0 0 0 0 8 3 0 0 4
566 241
590 241
590 169
597 169
2 7 5 0 0 0 0 4 9 0 0 4
427 176
426 176
426 241
424 241
3 0 15 0 0 0 0 8 0 0 35 3
512 250
487 250
487 302
3 0 15 0 0 0 0 9 0 0 35 3
370 250
340 250
340 302
4 3 15 0 0 8320 0 6 7 0 0 5
191 266
191 302
641 302
641 250
674 250
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
